// Serial Peripheral Interface virtual component

module

endmodule
