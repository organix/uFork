/*

Operation Encoding for ALU

*/

`ifndef _alu_ops_
`define _alu_ops_

`define NO_OP   (4'h0)
`define ADD_OP  (4'h1)
`define SUB_OP  (4'h2)
`define MUL_OP  (4'h3)
`define AND_OP  (4'h4)
`define XOR_OP  (4'h5)
`define OR_OP   (4'h6)
`define ROL_OP  (4'h7)

`endif
