/*
  Serial Peripheral Interface master virtual component

    +-----------------+
    | spi master      |
    |                 |
--->|i_spi_en   o_SCLK|--->
=8=>|i_data     o_MOSI|--->
<=8=|o_data     i_MISO|<---
<---|o_ready      o_SS|--->
    |                 |
 +->|i_clk            |
 |  +-----------------+

*/

module

endmodule
